`ifndef AXIMasterSlaveStream_v1_0_tb_include_vh_
`define AXIMasterSlaveStream_v1_0_tb_include_vh_

//Configuration current bd names
`define BD_NAME AXIMasterSlaveStreamIP_v1_0_bfm_1
`define BD_INST_NAME AXIMasterSlaveStreamIP_v1_0_bfm_1_i
`define BD_WRAPPER AXIMasterSlaveStreamIP_v1_0_bfm_1_wrapper

//Configuration address parameters
`endif
